module hello;
	initial begin
		$display("hello RISC-v");
		$finish;
	end
endmodule 
