module instruction_fetch_unit(
	input 
